module alu_8bit(
    input  wire [7:0] A,
    input  wire [7:0] B,
    input  wire [3:0] opcode,
    output reg  [7:0] result
);

    always @(*) begin
        case(opcode)
            4'b0000: result = A + B;           // ADD
            4'b0001: result = A - B;           // SUB
            4'b0010: result = A & B;           // AND
            4'b0011: result = A | B;           // OR
            4'b0100: result = A * B;           // MUL
            4'b0101: result = A ^ B;           // XOR
            4'b0110: result = A;               // PASS A
            4'b0111: result = B;               // PASS B
            4'b1000: result = A + 1;           // INC
            4'b1001: result = A - 1;           // DEC
            4'b1010: result = A << 1;          // SHIFT LEFT
            4'b1011: result = A >> 1;          // SHIFT RIGHT
            default: result = 8'h00;
        endcase
    end
endmodule
